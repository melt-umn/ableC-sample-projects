grammar bogus_table;

import edu:umn:cs:melt:ableC:host;

copper_mda testTablesTP(ablecParser) {
  bogus_table;
}

