grammar bogus_table_separator;

import edu:umn:cs:melt:ableC:host;

copper_mda testTablesTP(ablecParser) {
  bogus_table_separator;
}

