grammar artifact;

import edu:umn:cs:melt:ableC:drivers:compile;

construct ableC as
edu:umn:cs:melt:ableC:concretesyntax
translator using
  edu:umn:cs:melt:exts:ableC:run;
  edu:umn:cs:melt:exts:ableC:lvars;
  edu:umn:cs:melt:exts:ableC:templating;

  edu:umn:cs:melt:exts:ableC:run;
  edu:umn:cs:melt:exts:ableC:tensorAlgebra;

