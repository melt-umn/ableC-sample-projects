grammar bogus_scoped_table;

import edu:umn:cs:melt:ableC:host;

copper_mda testTablesTP(ablecParser) {
  bogus_scoped_table;
}

